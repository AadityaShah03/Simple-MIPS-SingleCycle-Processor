library verilog;
use verilog.vl_types.all;
entity mipsregisterfile_vlg_vec_tst is
end mipsregisterfile_vlg_vec_tst;
