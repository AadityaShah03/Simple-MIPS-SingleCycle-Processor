library verilog;
use verilog.vl_types.all;
entity nBitAddSub_vlg_vec_tst is
end nBitAddSub_vlg_vec_tst;
