library verilog;
use verilog.vl_types.all;
entity MIPS_ALU_8Bit_vlg_vec_tst is
end MIPS_ALU_8Bit_vlg_vec_tst;
