library verilog;
use verilog.vl_types.all;
entity decoder_3to8_vlg_vec_tst is
end decoder_3to8_vlg_vec_tst;
