library verilog;
use verilog.vl_types.all;
entity instrMem_vlg_vec_tst is
end instrMem_vlg_vec_tst;
