library verilog;
use verilog.vl_types.all;
entity nbit2to1mux_vlg_vec_tst is
end nbit2to1mux_vlg_vec_tst;
