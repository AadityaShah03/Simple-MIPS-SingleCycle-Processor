library verilog;
use verilog.vl_types.all;
entity Nbit_d_register_vlg_vec_tst is
end Nbit_d_register_vlg_vec_tst;
