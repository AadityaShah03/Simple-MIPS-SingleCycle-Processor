library verilog;
use verilog.vl_types.all;
entity DataMem_vlg_vec_tst is
end DataMem_vlg_vec_tst;
